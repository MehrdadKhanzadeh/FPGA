module adder (input [31:0] a, b, output reg [33:0] sum);

	assign sum = a + b;
	
endmodule	